* Created by KLayout

* cell Op8_18_rev1
* pin Bias
* pin Vdd
* pin OUT
* pin In+
* pin In1
* pin Vss
.SUBCKT Op8_18_rev1 11 14 15 19 22 26
* net 11 Bias
* net 14 Vdd
* net 15 OUT
* net 19 In+
* net 22 In1
* net 26 Vss
* device instance $1 r0 *1 42,79 NMOS
M$1 13 12 10 26 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $6 r0 *1 109,44 NMOS
M$6 1 2 26 26 NMOS L=5U W=20U AS=30P AD=30P PS=36U PD=36U
* device instance $8 r0 *1 95.5,44 NMOS
M$8 5 7 26 26 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $9 m90 *1 82,44 NMOS
M$9 6 7 26 26 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $10 m90 *1 32,49 NMOS
M$10 9 2 26 26 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $15 r0 *1 42,49 NMOS
M$15 10 2 26 26 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $20 r0 *1 93.5,69 NMOS
M$20 3 7 5 26 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $25 m90 *1 84,69 NMOS
M$25 7 7 6 26 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $30 m90 *1 138,44 NMOS
M$30 4 4 26 26 NMOS L=1U W=40U AS=50P AD=50P PS=60U PD=60U
* device instance $34 m90 *1 138,62 NMOS
M$34 8 8 4 26 NMOS L=1U W=40U AS=50P AD=50P PS=60U PD=60U
* device instance $38 m90 *1 32,79 NMOS
M$38 2 12 9 26 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $43 r0 *1 156.5,102.5 NMOS
M$43 15 27 15 26 NMOS L=1U W=100U AS=150P AD=150P PS=156U PD=156U
* device instance $45 r180 *1 145.5,104 NMOS
M$45 3 8 17 26 NMOS L=1U W=120U AS=160P AD=160P PS=168U PD=168U
* device instance $48 m90 *1 57,127.5 NMOS
M$48 20 19 13 26 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $53 r0 *1 67.5,127.5 NMOS
M$53 21 22 13 26 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $58 r0 *1 112.5,190.5 PMOS
M$58 17 11 14 14 PMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $59 m90 *1 28.5,187.5 PMOS
M$59 24 11 14 14 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $61 r0 *1 40,161 PMOS
M$61 12 11 25 14 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $66 m90 *1 133.5,152.5 PMOS
M$66 1 1 23 14 PMOS L=1U W=80U AS=100P AD=100P PS=110U PD=110U
* device instance $70 m90 *1 136,185.5 PMOS
M$70 23 23 14 14 PMOS L=1U W=80U AS=100P AD=100P PS=110U PD=110U
* device instance $74 r0 *1 41.5,187.5 PMOS
M$74 25 11 14 14 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $76 r0 *1 71.5,188 PMOS
M$76 21 11 14 14 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $78 r0 *1 91.5,188 PMOS
M$78 20 11 14 14 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $80 r0 *1 69,160.5 PMOS
M$80 7 11 21 14 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $85 m90 *1 30,161 PMOS
M$85 11 11 24 14 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $90 r0 *1 96,160.5 PMOS
M$90 18 11 20 14 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $95 r0 *1 149.5,165.5 PMOS
M$95 15 18 14 14 PMOS L=1U W=300U AS=360P AD=360P PS=372U PD=372U
* device instance $100 m90 *1 119.5,107.5 PMOS
M$100 3 1 18 14 PMOS L=1U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $105 r90 *1 78.5,103.5 HRES
R$105 12 2 17500 HRES
* device instance $106 r0 *1 254.75,59 CAP
C$106 15 3 9.49e-13 CAP
* device instance $108 m0 *1 254.75,172.5 CAP
C$108 15 18 9.49e-13 CAP
* device instance $112 r270 *1 37.5,103.5 HRES
R$112 26 11 350000 HRES
.ENDS Op8_18_rev1
