* Created by KLayout

* cell op8_18_v2_for_PTS06_LVS
* pin Bias
* pin OUT
* pin Vdd
* pin In+
* pin In1
* pin Vss
.SUBCKT op8_18_v2_for_PTS06_LVS 11 15 16 18 21 25
* net 11 Bias
* net 15 OUT
* net 16 Vdd
* net 18 In+
* net 21 In1
* net 25 Vss
* device instance $1 r0 *1 42,79 NMOS
M$1 13 12 8 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $6 m90 *1 73.5,44 NMOS
M$6 9 1 25 25 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $7 r0 *1 87.5,44 NMOS
M$7 10 1 25 25 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $8 m90 *1 84,69 NMOS
M$8 1 1 9 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $13 r0 *1 93.5,69 NMOS
M$13 5 1 10 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $18 m90 *1 32,49 NMOS
M$18 7 4 25 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $23 r0 *1 42,49 NMOS
M$23 8 4 25 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $28 m90 *1 145.5,59 NMOS
M$28 6 6 3 25 NMOS L=1U W=40U AS=50P AD=50P PS=60U PD=60U
* device instance $32 m90 *1 153,44 NMOS
M$32 3 3 25 25 NMOS L=1U W=40U AS=50P AD=50P PS=60U PD=60U
* device instance $36 m90 *1 32,79 NMOS
M$36 4 12 7 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $41 r0 *1 99.5,44 NMOS
M$41 2 4 25 25 NMOS L=5U W=60U AS=70P AD=70P PS=84U PD=84U
* device instance $47 r180 *1 161,100.5 NMOS
M$47 25 5 15 25 NMOS L=1U W=100U AS=150P AD=150P PS=156U PD=156U
* device instance $49 m90 *1 57,127.5 NMOS
M$49 19 18 13 25 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $54 r0 *1 67.5,127.5 NMOS
M$54 20 21 13 25 NMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $59 m90 *1 141.5,103.5 NMOS
M$59 17 6 5 25 NMOS L=1U W=120U AS=160P AD=160P PS=168U PD=168U
* device instance $62 m90 *1 122.5,107.5 PMOS
M$62 5 2 17 16 PMOS L=1U W=240U AS=280P AD=280P PS=294U PD=294U
* device instance $68 r0 *1 112.5,190.5 PMOS
M$68 6 11 16 16 PMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $69 m90 *1 28.5,187.5 PMOS
M$69 23 11 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $71 r0 *1 40,161 PMOS
M$71 12 11 24 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $76 m90 *1 133.5,152.5 PMOS
M$76 2 2 22 16 PMOS L=1U W=80U AS=100P AD=100P PS=110U PD=110U
* device instance $80 m90 *1 136,185.5 PMOS
M$80 22 22 16 16 PMOS L=1U W=80U AS=100P AD=100P PS=110U PD=110U
* device instance $84 r0 *1 71.5,188 PMOS
M$84 20 11 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $86 r0 *1 41.5,187.5 PMOS
M$86 24 11 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $88 r0 *1 91.5,188 PMOS
M$88 19 11 16 16 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $90 r0 *1 69,160.5 PMOS
M$90 1 11 20 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $95 m90 *1 30,161 PMOS
M$95 11 11 23 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $100 r0 *1 96,160.5 PMOS
M$100 17 11 19 16 PMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $105 r0 *1 149.5,165.5 PMOS
M$105 15 17 16 16 PMOS L=1U W=300U AS=360P AD=360P PS=372U PD=372U
* device instance $112 r270 *1 37.5,103.5 HRES
R$112 25 11 200000 HRES
* device instance $114 r90 *1 78.5,103.5 HRES
R$114 12 4 10000 HRES
* device instance $115 r0 *1 239.75,60.05 CAP
C$115 15 5 3.64e-13 CAP
* device instance $116 m0 *1 239.75,171.45 CAP
C$116 15 17 3.64e-13 CAP
.ENDS op8_18_v2_for_PTS06_LVS
